
module PS2 (
	clk_clk,
	reset_reset_n,
	ps2_0_external_interface_CLK,
	ps2_0_external_interface_DAT);	

	input		clk_clk;
	input		reset_reset_n;
	inout		ps2_0_external_interface_CLK;
	inout		ps2_0_external_interface_DAT;
endmodule
